---------------------------------------------------------------------------------
----! @file       ECC_MC_ROM.vhd
----! @brief      ECC Multiplier Scheduler ROM
----!
----! @author     Ahmed Ferozpuri
----! @copyright  Copyright (c) 2016 Cryptographic Engineering Research Group
----!             ECE Department, George Mason University Fairfax, VA, U.S.A.
----!             All rights Reserved.
---------------------------------------------------------------------------------
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
--
--entity ECC_MC_ROM is
	--port (
			--addr : in std_logic_vector (5 downto 0); -- address input
			--dout : out std_logic_vector (26 downto 0)); -- data output
--end ECC_MC_ROM;
 --
--architecture behave of ECC_MC_ROM is
 --
--type ECC_MC_ROMTABLE is array (0 to 41) of std_logic_vector (26 downto 0);
 ---- internal table
--constant romdata : ECC_MC_ROMTABLE := (
--"101010100000000000000000010",
--"000100000001000000000000101",
--"010010010000000000000000010",
--"001000100000000000000000010",
--"001100110000000000000000010",
--"000100010000000000000000010",
--"100101110111000000000000010",
--"101000101001000000000000010",
--"100110010111101101011010001",
--"100100111001000000000000010",
--"110010111011110101101001001",
--"101010101100000000000000010",
--"110011001011111010101010000",
--"011101111011111011001110000",
--"101111011101000000000000010",
--"100110011100010110111110001",
--"100001110111101010100101001",
--"101111011010000000000000010",
--"100010001000011010111001001",
--"100000011000000000000000010",
--"100101100110101001010101000",
--"101110011001101010101010000",
--"100110101001101110111011000",
--"101001010101101110111011000",
--"110001100111101110111011000",
--"110110111000111010101010000",
--"101011101010000000000000100",
--"101010101000000000000000100",
--"111010101010011111001100000",
--"110010011001000000000000100",
--"010111101100000000000000101",
--"100110010101000000000000101",
--"101010101001100011011101000",
--"011010101011000000000000101",
--"101010101010000000000000010",
--"101010100111000000000000010",
--"101110101010000000000000010",
--"001001011011000000000000010",
--"101110101011000000000000010",
--"001101101011000000000000010",
--"001010010010000000000000010",
--"001110010011000000000000010"
--);
 --
--begin
--
--process (addr)
--begin
	--dout <= romdata(to_integer(unsigned(addr)));
--end process;
 --
--end behave;

-------------------------------------------------------------------------------
--! @file       ECC_MC_ROM.vhd
--! @brief      ECC Multiplier Scheduler ROM
--!
--! @author     Ahmed Ferozpuri
--! @copyright  Copyright (c) 2016 Cryptographic Engineering Research Group
--!             ECE Department, George Mason University Fairfax, VA, U.S.A.
--!             All rights Reserved.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ECC_MC_ROM is
	port (
			addr : in std_logic_vector (6 downto 0); -- address input
			dout : out std_logic_vector (26 downto 0)); -- data output
end ECC_MC_ROM;
 
architecture behave of ECC_MC_ROM is
 
type ECC_MC_ROMTABLE is array (0 to 116) of std_logic_vector (26 downto 0);
 -- internal table
constant romdata : ECC_MC_ROMTABLE := (
"101000001010000000000000010", --0
"000100000001000000000000101", --1
"010010010000000000000000010", --2
"001000100000000000000000010", --3
"001100110000000000000000010", --4
"000111000000000000000000010", --5
"010001000011000000000000010", --6
"001100110011010001000100000", --7
"001100110011000000000000100", --8
"100100100010101100110010000", --9
"101110111011101010011001000", --10
"001100110011101110111001001", --11
"100110101001000000000000100", --12
"100100011001000000000000100", --13
"101010011001101110110011001", --14
"001010111011000000000000100", --15
"001010100010000000000000101", --16
"001100110011000000000000100", --17
"000100110001101110110010001", --18
"101110011011000100010001000", --19
"001110110011000000000000101", --20
"100101000100100001000111000", --21
"100010001000000000000000010", --22
"101001110111100010001001001", --23
"101101111010000000000000010", --24
"010101011001011110001010001", --25
"101000101010000000000000010", --26
"100101001001010101011010001", --27
"100101101001000000000000010", --28
"011000111011000000000000010", --29
"011101010111101101010101000", --30
"101110111011100110010110001", --31
"101010111010000000000000010", --32
"010110110101100110011001000", --33
"100010011001101110101010000", --34
"011001010110100010000101001", --35
"100001110111010110001011001", --36
"100010001000101010100101001", --37
"101010011010011001100110000", --38
"100011001000011010100110001", --39
"010001000011000000000000010", --40
"001100110011010001000100000", --41
"001100110011000000000000100", --42
"100100100010101100110010000", --43
"101110111011101010011001000", --44
"001100110011101110111001001", --45
"100110101001000000000000100", --46
"100100011001000000000000100", --47
"101010011001101110110011001", --48
"001010111011000000000000100", --49
"001010100010000000000000101", --50
"001100110011000000000000100", --51
"000100110001101110110010001", --52
"101110011011000100010001000", --53
"001110110011000000000000101", --54
"100101110111000101110100000", --55
"000100010001000000000000010", --56
"101001000100000100011001001", --57
"101101001010000000000000010", --58
"001000101001010000011010001", --59
"101001011010000000000000010", --60
"100101111001001000101010001", --61
"100100111001000000000000010", --62
"001101101011000000000000010", --63
"010000100100101100100010000", --64
"101110111011100110010011001", --65
"101010111010000000000000010", --66
"001010110010100110011001000", --67
"000110011001101110101010000", --68
"001100100011000100010010001", --69
"000101000100001000011011001", --70
"000100010001101010100010001", --71
"101010011010001100110011000", --72
"000111000001001110100011001", --73
"011101110110000000000000010", --74
"011001100110011101110111000", --75
"011001100110000000000000100", --76
"100101010101101101100101000", --77
"101110111011101010011001000", --78
"011001100110101110111001001", --79
"100110101001000000000000100", --80
"100110001001000000000000100", --81
"101010011001101110110110001", --82
"010110111011000000000000100", --83
"010110100101000000000000101", --84
"011001100110000000000000100", --85
"100001101000101110110101001", --86
"101110011011100010001000000", --87
"011010110110000000000000101", --88
"011011100110000000000000101", --89
"100111011101100011010111000", --90
"100010001000000000000000010", --91
"101001110111100010001001001", --92
"101101111010000000000000010", --93
"010101011001011110001010001", --94
"101000101010000000000000010", --95
"100111011001010101011010001", --96
"100101101001000000000000010", --97
"011000111011000000000000010", --98
"011101010111101101010101000", --99
"101110111011100110010110001", --100
"101010111010000000000000010", --101
"010110110101100110011001000", --102
"100010011001101110101010000", --103
"011001010110100010000101001", --104
"100001110111010110001011001", --105
"100010001000101010100101001", --106
"101010011010011001100110000", --107
"100011001000011010100110001", --108
"101010101010000000000000010", --109
"101010100111000000000000010", --110
"101110101010000000000000010", --111
"001001011011000000000000010", --112
"101110101011000000000000010", --113
"001101101011000000000000010", --114
"001010010010000000000000010", --115
"001110010011000000000000010"  --116
);
 
begin

process (addr)
begin
	dout <= romdata(to_integer(unsigned(addr)));
end process;
 
end behave;